library IEEE;
use IEEE.std_logic_1164.all;

package minesweeper_pkg is
    type natural_array is array(63 downto 0) of natural;
end package minesweeper_pkg;