library IEEE;
use IEEE.std_logic_1164.all;

package minesweeper_pkg is
    type number_array is array(63 downto 0) of std_logic_vector(3 downto 0);
end package minesweeper_pkg;